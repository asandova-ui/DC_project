//-------------------------------------------------------------------

//-------------------------------------------------------------------
`include "system.v"
`define SIMULATION

module tb();

//-- Registros con señales de entrada
reg clk;
reg resetb;
reg rxd;
wire txd;
integer k;
//-- Instanciamos 

SYSTEM sys1(	.clk(clk),		// Main clock input 25MHz
	.reset(~resetb),
	.rxd(rxd)
);

// Reloj periódico
always #5 clk=~clk;

//-- Proceso al inicio
initial begin
	//-- Fichero donde almacenar los resultados
	$dumpfile("tb.vcd");
	$dumpvars(0, tb);
		$dumpvars(0, tb.sys1.cpu.regs[11]);		
		$dumpvars(0, tb.sys1.cpu.regs[12]);		
		$dumpvars(0, tb.sys1.cpu.regs[13]);		
		$dumpvars(0, tb.sys1.cpu.regs[14]);		
		$dumpvars(0, tb.sys1.cpu.regs[15]);		

	resetb = 0; clk=0; rxd=1;

	#77		resetb=1;
	#10000  rxd=0;	//START
	
	#1560   rxd=1;
	#1560   rxd=0;
	#1560   rxd=0;
	#1560   rxd=0;

	#1560   rxd=0;
	#1560   rxd=0;
	#1560   rxd=1;
	#1560   rxd=0;

	#1560   rxd=1;	//STOP
	
	# 319 $display("FIN de la simulacion");
	//# 300000 $finish;
	# 1000 $finish;
end



endmodule


